







        















    









 







 



********************************        ****************************































































 




 










































  








 
 

  










  






 
 

  










  















           
















        
  







  






    











																																																																																																																						   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																									                           																																 			                                												      																																								    		    																			         									      									           																																																																																										    																																													                      																																																																																																																															           																																																																  				                                                    																																																																																																																										                                                                                							                                                                     																																																																																																																																																																																																																																																													                                																							    																																																																																																																																																																																																																																																																																																                                    								                     																																																																																																																																																																					  																													                                       																																																																																																																																																																																																																																											   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																							                   																																																																																																																																																																																																																																																																																																																																																																																																																																																																																					  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																															          																																																																																																																																																																																																							************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************                      ***********************************************************                                     *****************************         ************************************************************************************************************************************************************************************************************************************************************************************************************************************************************                                                                                                    ************************************************************************************************************  


 


 


 






 


 


 



























































































 

 



















































																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																														                  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																				      																																																																																																																																																																																																																																																																																																																																																																																																																																																																											      																																																																																																																																	                                ......................................................................................................................................................................................................................................................................................                                                                         .............................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................  ............................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                                                                                ......................................................................................................................................................................................................................................................................              ............................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                            